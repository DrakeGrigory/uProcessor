//ALU
`define ADD 3'd0
`define SUB 3'd1
`define AND 3'd2
`define OR  3'd3
`define XOR 3'd4
`define NOT 3'd5
`define LD  3'd6
